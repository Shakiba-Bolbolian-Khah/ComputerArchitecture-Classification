`timescale 1ns/1ns
module adder( input [13:0] op1, op2, output [13:0] result );
  assign result = op1 + op2;
endmodule
